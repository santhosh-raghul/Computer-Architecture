`include "fp-multiplier.v"

module top;

	reg [31:0]a, b;
	wire [31:0]out;

	m_fp_multiplier FP1 (a, b, out);

	initial
	begin

		a=32'b0_10001000_11101100000101000000100;	// 984.156494140625
		b=32'b0_10001011_01101110110100100101010;	// 5869.1455078125
		#5 $display("%b_%b_%b", out[31], out[30:23], out[22:0]);


		a=32'b1_10001011_00000100010111100100111;	// -4165.89404296875
		b=32'b0_10000110_00111000011000001110111;	// 156.18931579589844
		#5 $display("%b_%b_%b", out[31], out[30:23], out[22:0]);


		a=32'b1_10001100_10010101011110010100000;	// -12975.15625
		b=32'b1_10001110_01101111000011000110000;	// -46982.1875
		#5 $display("%b_%b_%b", out[31], out[30:23], out[22:0]);

	end

endmodule