`include "fp-adder.v"

module top;

	reg [31:0]a, b;
	wire [31:0]out;

	fp_adder FP1 (a, b, out);

	initial
begin

	// +ve +ve 
	a = 32'b0_10000000_11110000000000000000000;		// 3.875
	b = 32'b0_10000000_11000000000000000000000;		// 3.5
	// ==> 32'b0_10000001_11011000000000000000000  ans = 7.375

	
	// a = 32'b1_10000000_11000000000000000000000;		// 3.5
	// b = 32'b1_10000000_11000000000000000000000;		// 3.5
	
	// -ve -ve
	// a =	32'b1_10000010_00111000000000000000000;
	// b =	32'b1_10000010_00111000000000000000000;

	// a = 32'b0_10000010_00111000000000000000000;
	// b = 32'b0_10000000_11000000000000000000000;
	
	// infinity case
	// a = 32'b0_11111111_00000000000000000000000;
	// b = 32'b1_11111100_00000000000000000000000;

	// a = 32'b0_11111111_00000000000000000000000;
	// b = 32'b0_11111111_00000000000000000000000;

	// a = 32'b0_01111110_00100000000000000000000;
	// b = 32'b1_01111110_00100000000000000000000;

	// b = 32'b0_01111111_00000000000000000000000;
	// a = 32'h0000;
	// b = 32'h0000;

	#5 $display("ouS: %b %b %b", out[31], out[30:23], out[22:0]);
end

endmodule

// module top;

// 	reg [23:0]a;
// 	reg [4:0]s;
// 	wire [23:0]b;

// 	integer i;
// 	right_shift l(a,s,b);

// 	initial
// 	begin
// 		a = 24'b111111111111111111111111;
// 		for(i=0;i<32;i=i+1)
// 		begin
// 			s=i;
// 			#10 $display("%b %d %b",a,s,b);
// 		end
// 	end

// endmodule

// module top;

// 	reg [24:0]a;
// 	reg [4:0]s;
// 	wire [24:0]b,aw;

// 	integer i;
// 	left_shift l(aw,s,b);

// 	assign aw=a;
// 	initial
// 	begin
// 		a = 25'b1111111111111111111111111;
// 		for(i=0;i<32;i=i+1)
// 		begin
// 			s=i;
// 			#10 $display("%b %d %b",aw,s,b);
// 		end
// 	end

// endmodule